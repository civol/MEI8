library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity v95v95v58v840v58v58progv58v840v95e is
   port (
      addr: in std_logic_vector(7 downto 0);
      instr: out std_logic_vector(7 downto 0)
   );
end v95v95v58v840v58v58progv58v840v95e;

architecture v95v95v58v840v58v58progv58v840v95a of v95v95v58v840v58v58progv58v840v95e is

   type v58165 is array (0 to 255) of std_logic_vector(7 downto 0);
   constant content: v58165 := ( "00110110",
      "10101000",
      "10110100",
      "11111001",
      "10100101",
      "10110110",
      "11111001",
      "10101100",
      "10110110",
      "11111001",
      "10101100",
      "10110110",
      "11111001",
      "10101111",
      "10110110",
      "11111001",
      "10100001",
      "10110010",
      "11111001",
      "00000000",
      "00000000",
      "10100000",
      "10110010",
      "00000001",
      "10111000",
      "11111001",
      "01001001",
      "11101110",
      "00000000",
      "00000000",
      "10100101",
      "10111010",
      "00000010",
      "10100110",
      "01000010",
      "11111001",
      "00000011",
      "01010011",
      "01100011",
      "11111001",
      "00000100",
      "01011100",
      "01101100",
      "11111011",
      "00000101",
      "01110101",
      "10010101",
      "10000000",
      "11100010",
      "10010010",
      "10010000",
      "11010010",
      "10010000",
      "10010011",
      "11011010",
      "10010000",
      "10010100",
      "11001010",
      "10010000",
      "10010101",
      "10001101",
      "00101000",
      "10010000",
      "11110000",
      "10010000",
      "11110001",
      "10010000",
      "11110010",
      "10010000",
      "10111100",
      "11110100",
      "10010000",
      "11110011",
      "10010000",
      "11110110",
      "11111000",
      "10010000",
      "11111010",
      "10010000",
      "11111100",
      "11111110",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "00000000",
      "10100011",
      "11110111",
      "11111101",
      "00000000",
      "10101011",
      "10110100",
      "10011000",
      "11111111" );
begin
   instr <= content(to_integer(unsigned(addr)));

end v95v95v58v840v58v58progv58v840v95a;

